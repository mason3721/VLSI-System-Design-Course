`define CPU_CYCLE     9.8 // 100Mhz
`define MAX           1970000 // 3000000
