`define CPU_CYCLE     10.0 // 100Mhz
`define MAX           3000000 // 3000000
`define AXI_CYCLE     25.0 // 40Mhz
